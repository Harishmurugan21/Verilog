module buf_gate(input a,output y);
buf (y,a);
endmodule
