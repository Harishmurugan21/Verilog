module buf_if1 (input a,control,output y);
bufif1 (y,a,control);
endmodule
