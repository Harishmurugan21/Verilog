module parity_checker (input [4:0]a ,output even_parity);

assign even_parity =^a;
endmodule
          
