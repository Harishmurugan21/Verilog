
module and_gate(input a,b,output c);
//gate primitive
and(c,a,b);
endmodule

