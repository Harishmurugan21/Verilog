module mux_4to1_arrayindex (input [3:0]a,input [1:0]sel,output y);

assign y=a[sel];       //combining input lines into single array and 
		       //select the ouput based on 2 bit select line by index:
		       
		       
		 

endmodule


